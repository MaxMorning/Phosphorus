module ColorConverter (
    input wire[7:0] color256,

    output wire [7:0] r_value,
    output wire [7:0] g_value,
    output wire [7:0] b_value
);

    reg [23:0] color_24_bit;

    assign r_value = color_24_bit[23:16];
    assign g_value = color_24_bit[15:8];
    assign b_value = color_24_bit[7:0];

    always @(*) begin
        case (color256)
            0: color_24_bit = 24'hffffff;
            1: color_24_bit = 24'hffffcc;
            2: color_24_bit = 24'hffff99;
            3: color_24_bit = 24'hffff66;
            4: color_24_bit = 24'hffff33;
            5: color_24_bit = 24'hffff00;
            6: color_24_bit = 24'hffccff;
            7: color_24_bit = 24'hffcccc;
            8: color_24_bit = 24'hffcc99;
            9: color_24_bit = 24'hffcc66;
            10: color_24_bit = 24'hffcc33;
            11: color_24_bit = 24'hffcc00;
            12: color_24_bit = 24'hff99ff;
            13: color_24_bit = 24'hff99cc;
            14: color_24_bit = 24'hff9999;
            15: color_24_bit = 24'hff9966;
            16: color_24_bit = 24'hff9933;
            17: color_24_bit = 24'hff9900;
            18: color_24_bit = 24'hff66ff;
            19: color_24_bit = 24'hff66cc;
            20: color_24_bit = 24'hff6699;
            21: color_24_bit = 24'hff6666;
            22: color_24_bit = 24'hff6633;
            23: color_24_bit = 24'hff6600;
            24: color_24_bit = 24'hff33ff;
            25: color_24_bit = 24'hff33cc;
            26: color_24_bit = 24'hff3399;
            27: color_24_bit = 24'hff3366;
            28: color_24_bit = 24'hff3333;
            29: color_24_bit = 24'hff3300;
            30: color_24_bit = 24'hff00ff;
            31: color_24_bit = 24'hff00cc;
            32: color_24_bit = 24'hff0099;
            33: color_24_bit = 24'hff0066;
            34: color_24_bit = 24'hff0033;
            35: color_24_bit = 24'hff0000;
            36: color_24_bit = 24'hccffff;
            37: color_24_bit = 24'hccffcc;
            38: color_24_bit = 24'hccff99;
            39: color_24_bit = 24'hccff66;
            40: color_24_bit = 24'hccff33;
            41: color_24_bit = 24'hccff00;
            42: color_24_bit = 24'hccccff;
            43: color_24_bit = 24'hcccccc;
            44: color_24_bit = 24'hcccc99;
            45: color_24_bit = 24'hcccc66;
            46: color_24_bit = 24'hcccc33;
            47: color_24_bit = 24'hcccc00;
            48: color_24_bit = 24'hcc99ff;
            49: color_24_bit = 24'hcc99cc;
            50: color_24_bit = 24'hcc9999;
            51: color_24_bit = 24'hcc9966;
            52: color_24_bit = 24'hcc9933;
            53: color_24_bit = 24'hcc9900;
            54: color_24_bit = 24'hcc66ff;
            55: color_24_bit = 24'hcc66cc;
            56: color_24_bit = 24'hcc6699;
            57: color_24_bit = 24'hcc6666;
            58: color_24_bit = 24'hcc6633;
            59: color_24_bit = 24'hcc6600;
            60: color_24_bit = 24'hcc33ff;
            61: color_24_bit = 24'hcc33cc;
            62: color_24_bit = 24'hcc3399;
            63: color_24_bit = 24'hcc3366;
            64: color_24_bit = 24'hcc3333;
            65: color_24_bit = 24'hcc3300;
            66: color_24_bit = 24'hcc00ff;
            67: color_24_bit = 24'hcc00cc;
            68: color_24_bit = 24'hcc0099;
            69: color_24_bit = 24'hcc0066;
            70: color_24_bit = 24'hcc0033;
            71: color_24_bit = 24'hcc0000;
            72: color_24_bit = 24'h99ffff;
            73: color_24_bit = 24'h99ffcc;
            74: color_24_bit = 24'h99ff99;
            75: color_24_bit = 24'h99ff66;
            76: color_24_bit = 24'h99ff33;
            77: color_24_bit = 24'h99ff00;
            78: color_24_bit = 24'h99ccff;
            79: color_24_bit = 24'h99cccc;
            80: color_24_bit = 24'h99cc99;
            81: color_24_bit = 24'h99cc66;
            82: color_24_bit = 24'h99cc33;
            83: color_24_bit = 24'h99cc00;
            84: color_24_bit = 24'h9999ff;
            85: color_24_bit = 24'h9999cc;
            86: color_24_bit = 24'h999999;
            87: color_24_bit = 24'h999966;
            88: color_24_bit = 24'h999933;
            89: color_24_bit = 24'h999900;
            90: color_24_bit = 24'h9966ff;
            91: color_24_bit = 24'h9966cc;
            92: color_24_bit = 24'h996699;
            93: color_24_bit = 24'h996666;
            94: color_24_bit = 24'h996633;
            95: color_24_bit = 24'h996600;
            96: color_24_bit = 24'h9933ff;
            97: color_24_bit = 24'h9933cc;
            98: color_24_bit = 24'h993399;
            99: color_24_bit = 24'h993366;
            100: color_24_bit = 24'h993333;
            101: color_24_bit = 24'h993300;
            102: color_24_bit = 24'h9900ff;
            103: color_24_bit = 24'h9900cc;
            104: color_24_bit = 24'h990099;
            105: color_24_bit = 24'h990066;
            106: color_24_bit = 24'h990033;
            107: color_24_bit = 24'h990000;
            108: color_24_bit = 24'h66ffff;
            109: color_24_bit = 24'h66ffcc;
            110: color_24_bit = 24'h66ff99;
            111: color_24_bit = 24'h66ff66;
            112: color_24_bit = 24'h66ff33;
            113: color_24_bit = 24'h66ff00;
            114: color_24_bit = 24'h66ccff;
            115: color_24_bit = 24'h66cccc;
            116: color_24_bit = 24'h66cc99;
            117: color_24_bit = 24'h66cc66;
            118: color_24_bit = 24'h66cc33;
            119: color_24_bit = 24'h66cc00;
            120: color_24_bit = 24'h6699ff;
            121: color_24_bit = 24'h6699cc;
            122: color_24_bit = 24'h669999;
            123: color_24_bit = 24'h669966;
            124: color_24_bit = 24'h669933;
            125: color_24_bit = 24'h669900;
            126: color_24_bit = 24'h6666ff;
            127: color_24_bit = 24'h6666cc;
            128: color_24_bit = 24'h666699;
            129: color_24_bit = 24'h666666;
            130: color_24_bit = 24'h666633;
            131: color_24_bit = 24'h666600;
            132: color_24_bit = 24'h6633ff;
            133: color_24_bit = 24'h6633cc;
            134: color_24_bit = 24'h663399;
            135: color_24_bit = 24'h663366;
            136: color_24_bit = 24'h663333;
            137: color_24_bit = 24'h663300;
            138: color_24_bit = 24'h6600ff;
            139: color_24_bit = 24'h6600cc;
            140: color_24_bit = 24'h660099;
            141: color_24_bit = 24'h660066;
            142: color_24_bit = 24'h660033;
            143: color_24_bit = 24'h660000;
            144: color_24_bit = 24'h33ffff;
            145: color_24_bit = 24'h33ffcc;
            146: color_24_bit = 24'h33ff99;
            147: color_24_bit = 24'h33ff66;
            148: color_24_bit = 24'h33ff33;
            149: color_24_bit = 24'h33ff00;
            150: color_24_bit = 24'h33ccff;
            151: color_24_bit = 24'h33cccc;
            152: color_24_bit = 24'h33cc99;
            153: color_24_bit = 24'h33cc66;
            154: color_24_bit = 24'h33cc33;
            155: color_24_bit = 24'h33cc00;
            156: color_24_bit = 24'h3399ff;
            157: color_24_bit = 24'h3399cc;
            158: color_24_bit = 24'h339999;
            159: color_24_bit = 24'h339966;
            160: color_24_bit = 24'h339933;
            161: color_24_bit = 24'h339900;
            162: color_24_bit = 24'h3366ff;
            163: color_24_bit = 24'h3366cc;
            164: color_24_bit = 24'h336699;
            165: color_24_bit = 24'h336666;
            166: color_24_bit = 24'h336633;
            167: color_24_bit = 24'h336600;
            168: color_24_bit = 24'h3333ff;
            169: color_24_bit = 24'h3333cc;
            170: color_24_bit = 24'h333399;
            171: color_24_bit = 24'h333366;
            172: color_24_bit = 24'h333333;
            173: color_24_bit = 24'h333300;
            174: color_24_bit = 24'h3300ff;
            175: color_24_bit = 24'h3300cc;
            176: color_24_bit = 24'h330099;
            177: color_24_bit = 24'h330066;
            178: color_24_bit = 24'h330033;
            179: color_24_bit = 24'h330000;
            180: color_24_bit = 24'h00ffff;
            181: color_24_bit = 24'h00ffcc;
            182: color_24_bit = 24'h00ff99;
            183: color_24_bit = 24'h00ff66;
            184: color_24_bit = 24'h00ff33;
            185: color_24_bit = 24'h00ff00;
            186: color_24_bit = 24'h00ccff;
            187: color_24_bit = 24'h00cccc;
            188: color_24_bit = 24'h00cc99;
            189: color_24_bit = 24'h00cc66;
            190: color_24_bit = 24'h00cc33;
            191: color_24_bit = 24'h00cc00;
            192: color_24_bit = 24'h0099ff;
            193: color_24_bit = 24'h0099cc;
            194: color_24_bit = 24'h009999;
            195: color_24_bit = 24'h009966;
            196: color_24_bit = 24'h009933;
            197: color_24_bit = 24'h009900;
            198: color_24_bit = 24'h0066ff;
            199: color_24_bit = 24'h0066cc;
            200: color_24_bit = 24'h006699;
            201: color_24_bit = 24'h006666;
            202: color_24_bit = 24'h006633;
            203: color_24_bit = 24'h006600;
            204: color_24_bit = 24'h0033ff;
            205: color_24_bit = 24'h0033cc;
            206: color_24_bit = 24'h003399;
            207: color_24_bit = 24'h003366;
            208: color_24_bit = 24'h003333;
            209: color_24_bit = 24'h003300;
            210: color_24_bit = 24'h0000ff;
            211: color_24_bit = 24'h0000cc;
            212: color_24_bit = 24'h000099;
            213: color_24_bit = 24'h000066;
            214: color_24_bit = 24'h000033;
            215: color_24_bit = 24'hee0000;
            216: color_24_bit = 24'hdd0000;
            217: color_24_bit = 24'hbb0000;
            218: color_24_bit = 24'haa0000;
            219: color_24_bit = 24'h880000;
            220: color_24_bit = 24'h770000;
            221: color_24_bit = 24'h550000;
            222: color_24_bit = 24'h440000;
            223: color_24_bit = 24'h220000;
            224: color_24_bit = 24'h110000;
            225: color_24_bit = 24'h00ee00;
            226: color_24_bit = 24'h00dd00;
            227: color_24_bit = 24'h00bb00;
            228: color_24_bit = 24'h00aa00;
            229: color_24_bit = 24'h008800;
            230: color_24_bit = 24'h007700;
            231: color_24_bit = 24'h005500;
            232: color_24_bit = 24'h004400;
            233: color_24_bit = 24'h002200;
            234: color_24_bit = 24'h001100;
            235: color_24_bit = 24'h0000ee;
            236: color_24_bit = 24'h0000dd;
            237: color_24_bit = 24'h0000bb;
            238: color_24_bit = 24'h0000aa;
            239: color_24_bit = 24'h000088;
            240: color_24_bit = 24'h000077;
            241: color_24_bit = 24'h000055;
            242: color_24_bit = 24'h000044;
            243: color_24_bit = 24'h000022;
            244: color_24_bit = 24'h000011;
            245: color_24_bit = 24'heeeeee;
            246: color_24_bit = 24'hdddddd;
            247: color_24_bit = 24'hbbbbbb;
            248: color_24_bit = 24'haaaaaa;
            249: color_24_bit = 24'h888888;
            250: color_24_bit = 24'h777777;
            251: color_24_bit = 24'h555555;
            252: color_24_bit = 24'h444444;
            253: color_24_bit = 24'h222222;
            254: color_24_bit = 24'h111111;
            255: color_24_bit = 24'h000000;
            default:  color_24_bit = 24'heeeeee;
        endcase
    end

    
endmodule