module ColorConverter (
    input wire[7:0] color256,

    output wire [7:0] r_value,
    output wire [7:0] g_value,
    output wire [7:0] b_value
);

    reg [23:0] color_24_bit;

    assign r_value = color_24_bit[23:16];
    assign g_value = color_24_bit[15:8];
    assign b_value = color_24_bit[7:0];

    always @(*) begin
        case (color256)
            0: color_24_bit = 24'h000000;
            1: color_24_bit = 24'h800000;
            2: color_24_bit = 24'h008000;
            3: color_24_bit = 24'h808000;
            4: color_24_bit = 24'h000080;
            5: color_24_bit = 24'h800080;
            6: color_24_bit = 24'h008080;
            7: color_24_bit = 24'hc0c0c0;
            8: color_24_bit = 24'h808080;
            9: color_24_bit = 24'hff0000;
            10: color_24_bit = 24'h00ff00;
            11: color_24_bit = 24'hffff00;
            12: color_24_bit = 24'h0000ff;
            13: color_24_bit = 24'hff00ff;
            14: color_24_bit = 24'h00ffff;
            15: color_24_bit = 24'hffffff;
            16: color_24_bit = 24'h000000;
            17: color_24_bit = 24'h00005f;
            18: color_24_bit = 24'h000087;
            19: color_24_bit = 24'h0000af;
            20: color_24_bit = 24'h0000d7;
            21: color_24_bit = 24'h0000ff;
            22: color_24_bit = 24'h005f00;
            23: color_24_bit = 24'h005f5f;
            24: color_24_bit = 24'h005f87;
            25: color_24_bit = 24'h005faf;
            26: color_24_bit = 24'h005fd7;
            27: color_24_bit = 24'h005fff;
            28: color_24_bit = 24'h008700;
            29: color_24_bit = 24'h00875f;
            30: color_24_bit = 24'h008787;
            31: color_24_bit = 24'h0087af;
            32: color_24_bit = 24'h0087d7;
            33: color_24_bit = 24'h0087ff;
            34: color_24_bit = 24'h00af00;
            35: color_24_bit = 24'h00af5f;
            36: color_24_bit = 24'h00af87;
            37: color_24_bit = 24'h00afaf;
            38: color_24_bit = 24'h00afd7;
            39: color_24_bit = 24'h00afff;
            40: color_24_bit = 24'h00d700;
            41: color_24_bit = 24'h00d75f;
            42: color_24_bit = 24'h00d787;
            43: color_24_bit = 24'h00d7af;
            44: color_24_bit = 24'h00d7d7;
            45: color_24_bit = 24'h00d7ff;
            46: color_24_bit = 24'h00ff00;
            47: color_24_bit = 24'h00ff5f;
            48: color_24_bit = 24'h00ff87;
            49: color_24_bit = 24'h00ffaf;
            50: color_24_bit = 24'h00ffd7;
            51: color_24_bit = 24'h00ffff;
            52: color_24_bit = 24'h5f0000;
            53: color_24_bit = 24'h5f005f;
            54: color_24_bit = 24'h5f0087;
            55: color_24_bit = 24'h5f00af;
            56: color_24_bit = 24'h5f00d7;
            57: color_24_bit = 24'h5f00ff;
            58: color_24_bit = 24'h5f5f00;
            59: color_24_bit = 24'h5f5f5f;
            60: color_24_bit = 24'h5f5f87;
            61: color_24_bit = 24'h5f5faf;
            62: color_24_bit = 24'h5f5fd7;
            63: color_24_bit = 24'h5f5fff;
            64: color_24_bit = 24'h5f8700;
            65: color_24_bit = 24'h5f875f;
            66: color_24_bit = 24'h5f8787;
            67: color_24_bit = 24'h5f87af;
            68: color_24_bit = 24'h5f87d7;
            69: color_24_bit = 24'h5f87ff;
            70: color_24_bit = 24'h5faf00;
            71: color_24_bit = 24'h5faf5f;
            72: color_24_bit = 24'h5faf87;
            73: color_24_bit = 24'h5fafaf;
            74: color_24_bit = 24'h5fafd7;
            75: color_24_bit = 24'h5fafff;
            76: color_24_bit = 24'h5fd700;
            77: color_24_bit = 24'h5fd75f;
            78: color_24_bit = 24'h5fd787;
            79: color_24_bit = 24'h5fd7af;
            80: color_24_bit = 24'h5fd7d7;
            81: color_24_bit = 24'h5fd7ff;
            82: color_24_bit = 24'h5fff00;
            83: color_24_bit = 24'h5fff5f;
            84: color_24_bit = 24'h5fff87;
            85: color_24_bit = 24'h5fffaf;
            86: color_24_bit = 24'h5fffd7;
            87: color_24_bit = 24'h5fffff;
            88: color_24_bit = 24'h870000;
            89: color_24_bit = 24'h87005f;
            90: color_24_bit = 24'h870087;
            91: color_24_bit = 24'h8700af;
            92: color_24_bit = 24'h8700d7;
            93: color_24_bit = 24'h8700ff;
            94: color_24_bit = 24'h875f00;
            95: color_24_bit = 24'h875f5f;
            96: color_24_bit = 24'h875f87;
            97: color_24_bit = 24'h875faf;
            98: color_24_bit = 24'h875fd7;
            99: color_24_bit = 24'h875fff;
            100: color_24_bit = 24'h878700;
            101: color_24_bit = 24'h87875f;
            102: color_24_bit = 24'h878787;
            103: color_24_bit = 24'h8787af;
            104: color_24_bit = 24'h8787d7;
            105: color_24_bit = 24'h8787ff;
            106: color_24_bit = 24'h87af00;
            107: color_24_bit = 24'h87af5f;
            108: color_24_bit = 24'h87af87;
            109: color_24_bit = 24'h87afaf;
            110: color_24_bit = 24'h87afd7;
            111: color_24_bit = 24'h87afff;
            112: color_24_bit = 24'h87d700;
            113: color_24_bit = 24'h87d75f;
            114: color_24_bit = 24'h87d787;
            115: color_24_bit = 24'h87d7af;
            116: color_24_bit = 24'h87d7d7;
            117: color_24_bit = 24'h87d7ff;
            118: color_24_bit = 24'h87ff00;
            119: color_24_bit = 24'h87ff5f;
            120: color_24_bit = 24'h87ff87;
            121: color_24_bit = 24'h87ffaf;
            122: color_24_bit = 24'h87ffd7;
            123: color_24_bit = 24'h87ffff;
            124: color_24_bit = 24'haf0000;
            125: color_24_bit = 24'haf005f;
            126: color_24_bit = 24'haf0087;
            127: color_24_bit = 24'haf00af;
            128: color_24_bit = 24'haf00d7;
            129: color_24_bit = 24'haf00ff;
            130: color_24_bit = 24'haf5f00;
            131: color_24_bit = 24'haf5f5f;
            132: color_24_bit = 24'haf5f87;
            133: color_24_bit = 24'haf5faf;
            134: color_24_bit = 24'haf5fd7;
            135: color_24_bit = 24'haf5fff;
            136: color_24_bit = 24'haf8700;
            137: color_24_bit = 24'haf875f;
            138: color_24_bit = 24'haf8787;
            139: color_24_bit = 24'haf87af;
            140: color_24_bit = 24'haf87d7;
            141: color_24_bit = 24'haf87ff;
            142: color_24_bit = 24'hafaf00;
            143: color_24_bit = 24'hafaf5f;
            144: color_24_bit = 24'hafaf87;
            145: color_24_bit = 24'hafafaf;
            146: color_24_bit = 24'hafafd7;
            147: color_24_bit = 24'hafafff;
            148: color_24_bit = 24'hafd700;
            149: color_24_bit = 24'hafd75f;
            150: color_24_bit = 24'hafd787;
            151: color_24_bit = 24'hafd7af;
            152: color_24_bit = 24'hafd7d7;
            153: color_24_bit = 24'hafd7ff;
            154: color_24_bit = 24'hafff00;
            155: color_24_bit = 24'hafff5f;
            156: color_24_bit = 24'hafff87;
            157: color_24_bit = 24'hafffaf;
            158: color_24_bit = 24'hafffd7;
            159: color_24_bit = 24'hafffff;
            160: color_24_bit = 24'hd70000;
            161: color_24_bit = 24'hd7005f;
            162: color_24_bit = 24'hd70087;
            163: color_24_bit = 24'hd700af;
            164: color_24_bit = 24'hd700d7;
            165: color_24_bit = 24'hd700ff;
            166: color_24_bit = 24'hd75f00;
            167: color_24_bit = 24'hd75f5f;
            168: color_24_bit = 24'hd75f87;
            169: color_24_bit = 24'hd75faf;
            170: color_24_bit = 24'hd75fd7;
            171: color_24_bit = 24'hd75fff;
            172: color_24_bit = 24'hd78700;
            173: color_24_bit = 24'hd7875f;
            174: color_24_bit = 24'hd78787;
            175: color_24_bit = 24'hd787af;
            176: color_24_bit = 24'hd787d7;
            177: color_24_bit = 24'hd787ff;
            178: color_24_bit = 24'hd7af00;
            179: color_24_bit = 24'hd7af5f;
            180: color_24_bit = 24'hd7af87;
            181: color_24_bit = 24'hd7afaf;
            182: color_24_bit = 24'hd7afd7;
            183: color_24_bit = 24'hd7afff;
            184: color_24_bit = 24'hd7d700;
            185: color_24_bit = 24'hd7d75f;
            186: color_24_bit = 24'hd7d787;
            187: color_24_bit = 24'hd7d7af;
            188: color_24_bit = 24'hd7d7d7;
            189: color_24_bit = 24'hd7d7ff;
            190: color_24_bit = 24'hd7ff00;
            191: color_24_bit = 24'hd7ff5f;
            192: color_24_bit = 24'hd7ff87;
            193: color_24_bit = 24'hd7ffaf;
            194: color_24_bit = 24'hd7ffd7;
            195: color_24_bit = 24'hd7ffff;
            196: color_24_bit = 24'hff0000;
            197: color_24_bit = 24'hff005f;
            198: color_24_bit = 24'hff0087;
            199: color_24_bit = 24'hff00af;
            200: color_24_bit = 24'hff00d7;
            201: color_24_bit = 24'hff00ff;
            202: color_24_bit = 24'hff5f00;
            203: color_24_bit = 24'hff5f5f;
            204: color_24_bit = 24'hff5f87;
            205: color_24_bit = 24'hff5faf;
            206: color_24_bit = 24'hff5fd7;
            207: color_24_bit = 24'hff5fff;
            208: color_24_bit = 24'hff8700;
            209: color_24_bit = 24'hff875f;
            210: color_24_bit = 24'hff8787;
            211: color_24_bit = 24'hff87af;
            212: color_24_bit = 24'hff87d7;
            213: color_24_bit = 24'hff87ff;
            214: color_24_bit = 24'hffaf00;
            215: color_24_bit = 24'hffaf5f;
            216: color_24_bit = 24'hffaf87;
            217: color_24_bit = 24'hffafaf;
            218: color_24_bit = 24'hffafd7;
            219: color_24_bit = 24'hffafff;
            220: color_24_bit = 24'hffd700;
            221: color_24_bit = 24'hffd75f;
            222: color_24_bit = 24'hffd787;
            223: color_24_bit = 24'hffd7af;
            224: color_24_bit = 24'hffd7d7;
            225: color_24_bit = 24'hffd7ff;
            226: color_24_bit = 24'hffff00;
            227: color_24_bit = 24'hffff5f;
            228: color_24_bit = 24'hffff87;
            229: color_24_bit = 24'hffffaf;
            230: color_24_bit = 24'hffffd7;
            231: color_24_bit = 24'hffffff;
            232: color_24_bit = 24'h080808;
            233: color_24_bit = 24'h121212;
            234: color_24_bit = 24'h1c1c1c;
            235: color_24_bit = 24'h262626;
            236: color_24_bit = 24'h303030;
            237: color_24_bit = 24'h3a3a3a;
            238: color_24_bit = 24'h444444;
            239: color_24_bit = 24'h4e4e4e;
            240: color_24_bit = 24'h585858;
            241: color_24_bit = 24'h606060;
            242: color_24_bit = 24'h666666;
            243: color_24_bit = 24'h767676;
            244: color_24_bit = 24'h808080;
            245: color_24_bit = 24'h8a8a8a;
            246: color_24_bit = 24'h949494;
            247: color_24_bit = 24'h9e9e9e;
            248: color_24_bit = 24'ha8a8a8;
            249: color_24_bit = 24'hb2b2b2;
            250: color_24_bit = 24'hbcbcbc;
            251: color_24_bit = 24'hc6c6c6;
            252: color_24_bit = 24'hd0d0d0;
            253: color_24_bit = 24'hdadada;
            254: color_24_bit = 24'he4e4e4;
            default:  color_24_bit = 24'heeeeee;
        endcase
    end

    
endmodule